** Profile: "SCHEMATIC1-Reg. trans"  [ C:\Users\Sistemas Urban\Google Drive\Fiuba\Circuitos 2\Agosto 2018\C2_OBLIG3\cc-cc-SCHEMATIC1-Reg. trans.sim ] 

** Creating circuit file "cc-cc-SCHEMATIC1-Reg. trans.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1500us 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\cc-cc-SCHEMATIC1.net" 


.END
